`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/12/2024 12:29:23 PM
// Design Name: 
// Module Name: MUX4x1_testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MUX4x1_testbench();
//reg [0:3] in;
//reg [1:0] s;
//wire w1, w2, out;
//MUX4X1 DUT(in,s, out);
//   initial begin
//   in[0] = 4'b1; in[1] = 4'b0; in[2] = 4'b0; in[3] = 4'b0 ; s[0] = 2'b0; s[1] = 2'b0;
//   #100
   
//   in[0] = 4'b1; in[1] = 4'b0; in[2] = 4'b0; in[3] = 4'b0 ;  s[0] = 2'b0; s[1] = 2'b1;
// end
endmodule
